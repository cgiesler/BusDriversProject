`define MATMULA 32'h00000000
`define MATMULB 32'h00000100
`define MATMULC 32'h00000200
`define MATDIMM 32'h00000600
`define MATDIMN 32'h00000700
`define MATDIMP 32'h00000800
`define MATMULF 32'h00000A00
`define MAXPOLF 32'h00000C00