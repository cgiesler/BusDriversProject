//Version 0.1, Based off of UW-Madison ECE 552's
//cpu top level testbench
module cpu_top_tb();

logic clk, rst_n, nextTransaction, ack, en, go;
logic [1:0] Interrupt; //Not used for single
logic [31:0] memDataOut, memAddr; //Not used until DMA set up



wire [31:0] PC;
wire [31:0] Inst;           /* This should be the 15 bits of the FF that
                                  stores instructions fetched from instruction memory
                               */
wire        RegWrite;       /* Whether register file is being written to */
wire [4:0]  WriteRegister;  /* What register is written */
wire [31:0] WriteData;      /* Data */
wire        MemWrite;       /* Similar as above but for memory */
wire        MemRead;
wire [31:0] MemAddress;
wire [31:0] MemData;

wire        halt;         /* halt executed and in Memory or writeback stage */
        
integer     inst_count;
integer     cycle_count;

integer     trace_file;
integer     sim_log_file;



cpu_top DUT(.*);


   /* Setup */
   initial begin
      $display("Hello world...simulation starting");
      $display("See verilogsim.log and verilogsim.trace for output");
      inst_count = 0;
      trace_file = $fopen("verilogsim.trace");
      sim_log_file = $fopen("verilogsim.log");
      
   end


  /* Clock and Reset */
// Clock period is 100 time units, and reset length
// to 201 time units (two rising edges of clock).

   initial begin
      $dumpvars;
      cycle_count = 0;
	  Interrupt = 2'b00;
      rst_n = 0; /* Intial reset state */
	  go = 0;
      clk = 1;
      #201 rst_n = 1; // delay until slightly after two clock periods
	  go = 1;
    end

    always #50 begin   // delay 1/2 clock period each time thru loop
      clk = ~clk;
    end
	
    always @(posedge clk) begin
    	cycle_count = cycle_count + 1;
	if (cycle_count > 100000) begin
		$display("hmm....more than 100000 cycles of simulation...error?\n");
		$finish;
	end
    end


/* Stats */
always @ (posedge clk) begin
	if (rst_n) begin
        	if (halt || RegWrite || MemWrite) begin
            	inst_count = inst_count + 1;
         	end
         	$fdisplay(sim_log_file, "SIMLOG:: Cycle %d PC: %8x I: %8x R: %d %3d %8x M: %d %d %8x %8x",
                cycle_count,
                PC,
                Inst,
                RegWrite,
                WriteRegister,
                WriteData,
                MemRead,
                MemWrite,
                MemAddress,
                MemData);
		if (RegWrite) begin
        	if (MemRead) begin
               	// ld
               	$fdisplay(trace_file,"INUM: %8d PC: 0x%04x REG: %d VALUE: 0x%04x ADDR: 0x%04x",
                         (inst_count-1),
                        PC,
                        WriteRegister,
                        WriteData,
                        MemAddress);
            	end else begin
               	$fdisplay(trace_file,"INUM: %8d PC: 0x%04x REG: %d VALUE: 0x%04x",
                         (inst_count-1),
                        PC,
                        WriteRegister,
                        WriteData );
            	end
		end else if (halt) begin
        	$fdisplay(sim_log_file, "SIMLOG:: Processor halted\n");
           	$fdisplay(sim_log_file, "SIMLOG:: sim_cycles %d\n", cycle_count);
           	$fdisplay(sim_log_file, "SIMLOG:: inst_count %d\n", inst_count);
           	$fdisplay(trace_file, "INUM: %8d PC: 0x%04x",
                      (inst_count-1),
                      PC );

           	$fclose(trace_file);
           	$fclose(sim_log_file);
            
           	$finish;
         end else begin
            	if (MemWrite) begin
               		// st
               		$fdisplay(trace_file,"INUM: %8d PC: 0x%04x ADDR: 0x%04x VALUE: 0x%04x",
                        (inst_count-1),
                        PC,
                        MemAddress,
                        MemData);
            	end else begin
            		// conditional branch or NOP
               		// Need better checking in pipelined testbench
               		inst_count = inst_count + 1;
               		$fdisplay(trace_file, "INUM: %8d PC: 0x%04x",
                         (inst_count-1),
                         PC );
            	end
		end 
	end      
end


   /* Assign internal signals to top level wires
      The internal module names and signal names will vary depending
      on your naming convention and your design */

   // Edit the example below. You must change the signal
   // names on the right hand side
    
//   assign PC = DUT.fetch0.pcCurrent; //You won't need this because it's part of the main cpu interface
   //assign Inst = DUT.fetch0.instr;
   assign Inst = DUT.inst;

   //assign RegWrite = DUT.decode0.regFile0.write;
   assign RegWrite = DUT.W_wEn;
   // Is memory being read, one bit signal (1 means yes, 0 means no)
   
   //assign WriteRegister = DUT.decode0.regFile0.writeregsel;
   assign WriteRegister = DUT.W_wReg;
   // The name of the register being written to. (4 bit signal)

   //assign WriteData = DUT.decode0.regFile0.writedata;
   assign WriteData = DUT.W_wData;
   // Data being written to the register. (16 bits)
   
   //assign MemRead =  DUT.memory0.memRead;
   assign MemRead =  DUT.M_memrd;
   // Is memory being read, one bit signal (1 means yes, 0 means no)
   
   //assign MemWrite = (DUT.memory0.memReadorWrite & DUT.memory0.memWrite);
   assign MemWrite = DUT.M_memwr;
   // Is memory being written to (1 bit signal)
   
   //assign MemAddress = DUT.memory0.aluResult;
   assign MemAddress = DUT.M_addrOut;
   // Address to access memory with (for both reads and writes to memory, 16 bits)
   
   //assign MemData = DUT.memory0.writeData;
   assign MemData = DUT.M_Reg1Out;
   // Data to be written to memory for memory writes (16 bits)
   
//   assign halt = DUT.memory0.halt; //You won't need this because it's part of the main cpu interface
   // Is processor halted (1 bit signal)
   
   /* Add anything else you want here */


endmodule

